// ============================================================================
// DE10-Lite Top Level Module
// ============================================================================

`define ENABLE_ADC_CLOCK
`define ENABLE_CLOCK1
`define ENABLE_CLOCK2
`define ENABLE_SDRAM
`define ENABLE_HEX0
`define ENABLE_HEX1
`define ENABLE_HEX2
`define ENABLE_HEX3
`define ENABLE_HEX4
`define ENABLE_HEX5
`define ENABLE_KEY
`define ENABLE_LED
`define ENABLE_SW
`define ENABLE_VGA
`define ENABLE_ACCELEROMETER
`define ENABLE_ARDUINO
`define ENABLE_GPIO

module DE10_LITE_Golden_Top(

	//////////// ADC CLOCK: 3.3-V LVTTL //////////
`ifdef ENABLE_ADC_CLOCK
	input 		          		ADC_CLK_10,
`endif
	//////////// CLOCK 1: 3.3-V LVTTL //////////
`ifdef ENABLE_CLOCK1
	input 		          		MAX10_CLK1_50,
`endif
	//////////// CLOCK 2: 3.3-V LVTTL //////////
`ifdef ENABLE_CLOCK2
	input 		          		MAX10_CLK2_50,
`endif

	//////////// SDRAM: 3.3-V LVTTL //////////
`ifdef ENABLE_SDRAM
	output		    [12:0]		DRAM_ADDR,
	output		     [1:0]		DRAM_BA,
	output		          		DRAM_CAS_N,
	output		          		DRAM_CKE,
	output		          		DRAM_CLK,
	output		          		DRAM_CS_N,
	inout 		    [15:0]		DRAM_DQ,
	output		          		DRAM_LDQM,
	output		          		DRAM_RAS_N,
	output		          		DRAM_UDQM,
	output		          		DRAM_WE_N,
`endif

	//////////// SEG7: 3.3-V LVTTL //////////
`ifdef ENABLE_HEX0
	output		     [7:0]		HEX0,
`endif
`ifdef ENABLE_HEX1
	output		     [7:0]		HEX1,
`endif
`ifdef ENABLE_HEX2
	output		     [7:0]		HEX2,
`endif
`ifdef ENABLE_HEX3
	output		     [7:0]		HEX3,
`endif
`ifdef ENABLE_HEX4
	output		     [7:0]		HEX4,
`endif
`ifdef ENABLE_HEX5
	output		     [7:0]		HEX5,
`endif

	//////////// KEY: 3.3 V SCHMITT TRIGGER //////////
`ifdef ENABLE_KEY
	input 		     [1:0]		KEY,
`endif

	//////////// LED: 3.3-V LVTTL //////////
`ifdef ENABLE_LED
	output		     [9:0]		LEDR,
`endif

	//////////// SW: 3.3-V LVTTL //////////
`ifdef ENABLE_SW
	input 		     [9:0]		SW,
`endif

	//////////// VGA: 3.3-V LVTTL //////////
`ifdef ENABLE_VGA
	output		     [3:0]		VGA_B,
	output		     [3:0]		VGA_G,
	output		          		VGA_HS,
	output		     [3:0]		VGA_R,
	output		          		VGA_VS,
`endif

	//////////// Accelerometer: 3.3-V LVTTL //////////
`ifdef ENABLE_ACCELEROMETER
	output		          		GSENSOR_CS_N,
	input 		     [2:1]		GSENSOR_INT,
	output		          		GSENSOR_SCLK,
	inout 		          		GSENSOR_SDI,
	inout 		          		GSENSOR_SDO,
`endif

	//////////// Arduino: 3.3-V LVTTL //////////
`ifdef ENABLE_ARDUINO
	inout 		    [15:0]		ARDUINO_IO,
	inout 		          		ARDUINO_RESET_N,
`endif

	//////////// GPIO, GPIO connect to GPIO Default: 3.3-V LVTTL //////////
`ifdef ENABLE_GPIO
	inout 		    [35:0]		GPIO
`endif
);



//=======================================================
//  REG/WIRE declarations
//=======================================================




//=======================================================
//  Structural coding
//=======================================================

	wire [6:0] hex0_seg, hex1_seg, hex2_seg, hex3_seg;
	wire [9:0] led_status;
	
	// Instantiate stopwatch module
	stopwatch_top u_stopwatch (
		.CLOCK_50(MAX10_CLK1_50),
		.KEY(KEY[1:0]),
		.HEX0(hex0_seg),
		.HEX1(hex1_seg),
		.HEX2(hex2_seg),
		.HEX3(hex3_seg),
		.LEDR(led_status)
	);
	
	// Connect 7-bit segment output to 8-bit HEX outputs (add decimal point)
	assign HEX0 = {1'b1, hex0_seg};  // Active-low, so 1 = off
	assign HEX1 = {1'b1, hex1_seg};
	assign HEX2 = {1'b1, hex2_seg};
	assign HEX3 = {1'b1, hex3_seg};
	assign HEX4 = 8'b11111111;       // Turn off HEX4
	assign HEX5 = 8'b11111111;       // Turn off HEX5

//=======================================================
//  Default assignments for unused outputs
//=======================================================

`ifdef ENABLE_LED
	// Connect LED status from stopwatch module
	assign LEDR = led_status;
`endif

`ifdef ENABLE_SDRAM
	// SDRAM - set to safe inactive state
	assign DRAM_ADDR  = 13'b0;
	assign DRAM_BA    = 2'b0;
	assign DRAM_CAS_N = 1'b1;       // Active-low, so 1 = inactive
	assign DRAM_CKE   = 1'b0;       // Clock enable off
	assign DRAM_CLK   = 1'b0;
	assign DRAM_CS_N  = 1'b1;       // Active-low, so 1 = deselected
	assign DRAM_LDQM  = 1'b1;       // Mask data
	assign DRAM_RAS_N = 1'b1;       // Active-low, so 1 = inactive
	assign DRAM_UDQM  = 1'b1;       // Mask data
	assign DRAM_WE_N  = 1'b1;       // Active-low, so 1 = no write
	// DRAM_DQ is inout - set to high-impedance
	assign DRAM_DQ    = 16'bz;
`endif

`ifdef ENABLE_VGA
	// VGA - blank screen (active video = 0)
	assign VGA_R  = 4'b0;
	assign VGA_G  = 4'b0;
	assign VGA_B  = 4'b0;
	assign VGA_HS = 1'b1;           // Sync signals idle high
	assign VGA_VS = 1'b1;
`endif

`ifdef ENABLE_ACCELEROMETER
	// Accelerometer - inactive state
	assign GSENSOR_CS_N  = 1'b1;    // Active-low, so 1 = deselected
	assign GSENSOR_SCLK  = 1'b0;    // Clock idle low
	// Bidirectional pins set to high-impedance
	assign GSENSOR_SDI   = 1'bz;
	assign GSENSOR_SDO   = 1'bz;
`endif

`ifdef ENABLE_ARDUINO
	// Arduino header - high-impedance (allow external use)
	assign ARDUINO_IO      = 16'bz;
	assign ARDUINO_RESET_N = 1'bz;
`endif

`ifdef ENABLE_GPIO
	// GPIO - high-impedance (allow external use)
	assign GPIO = 36'bz;
`endif

endmodule
